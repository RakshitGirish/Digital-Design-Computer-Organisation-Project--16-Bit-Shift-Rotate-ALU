module sll(input wire [15:0] i, input wire [3:0] shift_by, output wire [15:0] o);
    mux16 by15( { i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0] }, shift_by, o[15]);
	mux16 by14( { i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0 }, shift_by, o[14]);
    mux16 by13( { i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0 }, shift_by, o[13]);
    mux16 by12( { i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0 }, shift_by, o[12]);
    mux16 by11( { i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[11]);
    mux16 by10( { i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[10]);
    mux16 by9( { i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[9]);
    mux16 by8( { i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[8]);
    mux16 by7( { i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[7]);
    mux16 by6( { i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[6]);
    mux16 by5( { i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[5]);
    mux16 by4( { i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[4]);
    mux16 by3( { i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[3]);
    mux16 by2( { i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[2]);
    mux16 by1( { i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[1]);
    mux16 by0( { i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[0]);
endmodule

module srl(input wire [15:0] i, input wire [3:0] shift_by, output wire [15:0] o);
    mux16 by0( { i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15] }, shift_by, o[0]);
    mux16 by1( { i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0 }, shift_by, o[1]);
    mux16 by2( { i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0 }, shift_by, o[2]);
    mux16 by3( { i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0 }, shift_by, o[3]);
    mux16 by4( { i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[4]);
    mux16 by5( { i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[5]);
    mux16 by6( { i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[6]);
    mux16 by7( { i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[7]);
    mux16 by8( { i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[8]);
    mux16 by9( { i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[9]);
    mux16 by10( { i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[10]);
    mux16 by11( { i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[11]);
    mux16 by12( { i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[12]);
    mux16 by13( { i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[13]);
    mux16 by14( { i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[14]);
    mux16 by15( { i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift_by, o[15]);
endmodule

module rr(input wire [15:0] i, input wire [3:0] shift_by, output wire [15:0] o);
    mux16 by0( { i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15] }, shift_by, o[0]);
    mux16 by1( { i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0] }, shift_by, o[1]);
    mux16 by2( { i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1] }, shift_by, o[2]);
    mux16 by3( { i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2] }, shift_by, o[3]);
    mux16 by4( { i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3] }, shift_by, o[4]);
    mux16 by5( { i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4] }, shift_by, o[5]);
    mux16 by6( { i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5] }, shift_by, o[6]);
    mux16 by7( { i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6] }, shift_by, o[7]);
    mux16 by8( { i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7] }, shift_by, o[8]);
    mux16 by9( { i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8] }, shift_by, o[9]);
    mux16 by10( { i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8],i[9] }, shift_by, o[10]);
    mux16 by11( { i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10] }, shift_by, o[11]);
    mux16 by12( { i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11] }, shift_by, o[12]);
    mux16 by13( { i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12] }, shift_by, o[13]);
    mux16 by14( { i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13] }, shift_by, o[14]);
    mux16 by15( { i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14] }, shift_by, o[15]);
endmodule

module rl(input wire [15:0] i, input wire [3:0] shift_by, output wire [15:0] o);
    mux16 by15( { i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0] }, shift_by, o[15]);
    mux16 by14( { i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15]}, shift_by, o[14]);
    mux16 by13( { i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14] }, shift_by, o[13]);
    mux16 by12( { i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13] }, shift_by, o[12]);
    mux16 by11( { i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12] }, shift_by, o[11]);
    mux16 by10( { i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11] }, shift_by, o[10]);
    mux16 by9( { i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10] }, shift_by, o[9]);
    mux16 by8( { i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9] }, shift_by, o[8]);
    mux16 by7( { i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8] }, shift_by, o[7]);
    mux16 by6( { i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7] }, shift_by, o[6]);
    mux16 by5( { i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6] }, shift_by, o[5]);
    mux16 by4( { i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5] }, shift_by, o[4]);
    mux16 by3( { i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4] }, shift_by, o[3]);
    mux16 by2( { i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3] }, shift_by, o[2]);
    mux16 by1( { i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2] }, shift_by, o[1]);
    mux16 by0( { i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1] }, shift_by, o[0]);
endmodule

module alu (input wire [1:0] choice, input wire [15:0] i0, input wire [3:0] shift_by,output wire [15:0] o);
	wire [15:0] sll_op, srl_op, rr_op, rl_op;

    sll shift_left(i0, shift_by, sll_op);    
    rl rotate_left(i0, shift_by, rl_op);     
    srl shift_right(i0, shift_by, srl_op);   
    rr rotate_right(i0, shift_by, rr_op);    

    assign o = (choice[1] == 1'b0) ? ((choice[0] == 1'b0) ? sll_op : rl_op) : ((choice[0] == 1'b0) ? srl_op : rr_op);
endmodule
